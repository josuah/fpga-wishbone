module wbs_nvic #(
) (
);

endmodule
