interface iWishboneBus ( input logic clk, rst);
	iWishbone.controller wbc;
	iWishbone.peripheral wbp;
endinterface
